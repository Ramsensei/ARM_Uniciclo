module decoder(input logic [1:0] Op,
					input logic [5:0] Funct,
					input logic [3:0] Rd,
					output logic [1:0] FlagW,
					output logic PCS, RegW, MemW,
					output logic MemtoReg, ALUSrc,
					output logic [1:0] ImmSrc, RegSrc, ALUControl,
					output logic cs);
					
logic [9:0] controls;
logic Branch, ALUOp;
// Main Decoder
always_comb
casex(Op)
		// Data-processing immediate
		2'b00: if (Funct[5]) controls = 11'b00001010010;
		// Data-processing register
		else controls = 11'b00000010010;
		// LDR
		2'b01: if (Funct[0]) controls = 11'b00011110000;
		// STR
		else controls = 11'b10011101000;
		// B
		2'b10: controls = 11'b01101000100;
		// Unimplemented
		2'b11: controls = 11'b00000000001;
		default: controls = 11'bx;
endcase

assign {RegSrc, ImmSrc, ALUSrc, MemtoReg,
RegW, MemW, Branch, ALUOp, cs} = controls;

// ALU Decoder
always_comb
if (ALUOp) begin // which DP Instr?
case(Funct[4:1])
		4'b0100: ALUControl = 2'b00; // ADD
		4'b0010: ALUControl = 2'b01; // SUB
		4'b0000: ALUControl = 2'b10; // AND
		4'b1100: ALUControl = 2'b11; // ORR
		default: ALUControl = 2'bx;  // unimplemented
endcase

// update flags if S bit is set (C & V only for arith)
FlagW[1] = Funct[0];
FlagW[0] = Funct[0] &
	(ALUControl == 2'b00 | ALUControl == 2'b01);
end else begin
	ALUControl = 2'b00; // add for non-DP instructions
	FlagW = 2'b00; // don't update Flags
end
// PC Logic
	assign PCS = ((Rd == 4'b1111) & RegW) | Branch;
endmodule